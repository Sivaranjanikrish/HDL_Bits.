//Build a circuit with no inputs and one output that outputs a constant 
module constant0(out);
  output out;
	assign out=1'b0;
endmodule
